parameter KYBER_K = 256;
parameter KYBER_N = 3;
parameter KYBER_Q = 3329;
parameter KYBER_ETA = 2;
parameter KYBER_DU = 10;
parameter KYBER_DV = 4;
parameter KYBER_R_WIDTH = 12;


// HASH
parameter SHAKE_RATE = 1344;
parameter SHAKE_CAPACITY = 256;
parameter SHAKE_DOMAIN_SEPAROATOR = 8'h1F
