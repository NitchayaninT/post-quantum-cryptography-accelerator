`timescale 1ns/1ps
`include "params.vh"

module decode_pk_tb;

endmodule
