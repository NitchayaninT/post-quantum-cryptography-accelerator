// Kyber `define default we use Kyber-768
`define KYBER_K 3
`define KYBER_N 256
`define KYBER_Q 3329
`define KYBER_ETA 2
`define KYBER_DU 10
`define KYBER_DV 4
`define KYBER_R_WIDTH 12
`define KYBER_ARITH_W 16
`define KYBER_SPOLY_WIDTH 3

// HASH
`define SHAKE_RATE 1344
`define SHAKE_CAPACITY 256
`define SHAKE_DOMAIN_SEPAROATOR 8'h1F

`define DELAY 10
